library ieee;
use ieee.std_logic_1164.all;

entity g14_test is
port();
end g14_test;

architecture imp for g14_test is
--bla bla
begin
-- more bla bla
end imp;
